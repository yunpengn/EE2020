`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Niu Yunpeng
//////////////////////////////////////////////////////////////////////////////////

module my_dff(input CLOCK, input D, output reg OUT);
    always @(posedge CLOCK) begin
        OUT <= D;
    end
endmodule
